module fetch(clk, reset, new_addr, new_addr_valid, dram_en, dram_rdwr, dram_data, dram_addr, dram_valid);

endmodule
